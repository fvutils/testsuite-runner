/****************************************************************************
 * vlog_sim_smoke_tb.sv
 ****************************************************************************/

/**
 * Module: vlog_sim_smoke_tb
 * 
 * TODO: Add module documentation
 */
module vlog_sim_smoke_tb(input clk);

    initial begin
        $display("Hello World");
    end


endmodule


